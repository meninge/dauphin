LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
USE ieee.std_logic_unsigned.all;
Library UNISIM;
use UNISIM.vcomponents.all;
library UNIMACRO;
use unimacro.Vcomponents.all;

use iEEE.numeric_std.all;

-- entity declaration for your testbench.Dont declare any ports here
ENTITY test_1neuron_fsm IS 
	END test_1neuron_fsm;

ARCHITECTURE behavior OF test_1neuron_fsm IS
	-- add component under test
	component fsm
		generic ( NB_NEURONS : natural);
		port (
			     reset         : in  std_logic;
			     clk           : in  std_logic;
			     -- Control signals
			     ctrl_we_mode    : out  std_logic;
			     ctrl_we_shift   : out  std_logic;
			     ctrl_we_valid   : out  std_logic;
			     ctrl_accu_clear : out  std_logic;
			     ctrl_accu_add   : out  std_logic;
			     ctrl_shift_en   : out  std_logic;
			     ctrl_shift_copy : out  std_logic;
			     -- Address used for Read and Write
			     addr            : out  std_logic_vector(9 downto 0);
			     -- Ports for Write Enable
			     n0_we_prev         : out  std_logic;
			     nN_we_next         : in std_logic;
			     -- Sensors, for synchronization with the controller
			     sensor_shift    : in std_logic;
			     sensor_copy     : in std_logic;
			     sensor_we_mode  : in std_logic;
			     sensor_we_shift : in std_logic;
			     sensor_we_valid : in std_logic;

			     -- inputs
			     fsm_mode	: in std_logic;
			     -- in FIFO
			     cnt_fifo_in : in std_logic_vector(15 downto 0);
			     ack_fifo_in : out std_logic;
			     -- out FIFO
			     cnt_fifo_out  : in std_logic_vector(15 downto 0);
			     ack_fifo_out  : out std_logic
		     );
	end component;
	component neuron
		port(
			clk             : in  std_logic;
			-- Control signals
			ctrl_we_mode    : in  std_logic;
			ctrl_we_shift   : in  std_logic;
			ctrl_we_valid   : in  std_logic;
			ctrl_accu_clear : in  std_logic;
			ctrl_accu_add   : in  std_logic;
			ctrl_shift_en   : in  std_logic;
			ctrl_shift_copy : in  std_logic;
			-- Address used for Read and Write
			addr            : in  std_logic_vector(9 downto 0);
			-- Ports for Write Enable
			we_prev         : in  std_logic;
			we_next         : out std_logic;
			write_data      : in  std_logic_vector(15 downto 0);
			-- Data input, 2 bits
			data_in         : in  std_logic_vector(15 downto 0);
			-- Scan chain to extract values
			sh_data_in      : in  std_logic_vector(31 downto 0);
			sh_data_out     : out std_logic_vector(31 downto 0);
			-- Sensors, for synchronization with the controller
			sensor_shift    : out std_logic;
			sensor_copy     : out std_logic;
			sensor_we_mode  : out std_logic;
			sensor_we_shift : out std_logic;
			sensor_we_valid : out std_logic

		    );
	end component;
	

	signal clk           :   std_logic := '0';
	signal reset         :   std_logic := '0';
	-- Control signals
	signal ctrl_we_mode    :   std_logic := '0';
	signal ctrl_we_shift   :   std_logic := '0';
	signal ctrl_we_valid   :   std_logic := '0';
	signal ctrl_accu_clear :   std_logic := '0';
	signal ctrl_accu_add   :   std_logic := '0';
	signal ctrl_shift_en   :   std_logic := '0';
	signal ctrl_shift_copy :   std_logic := '0';
	-- Address used for Read and Write
	signal addr            :   std_logic_vector(9 downto 0);
	-- Ports for Write Enable
	signal n0_we_prev      :   std_logic := '0';
	signal nN_we_next      :  std_logic := '0';
	-- data weight
	signal write_data   :  std_logic_vector(15 downto 0);
	-- Data input, 2 bits
	signal data_in         : std_logic_vector(15 downto 0);
	-- Scan chain to extract values
	signal sh_data_in      : std_logic_vector(31 downto 0);
	signal sh_data_out     : std_logic_vector(31 downto 0);
	-- Sensors, for synchronization with the controller
	signal sensor_shift    :  std_logic := '0';
	signal sensor_copy     :  std_logic := '0';
	signal sensor_we_mode  :  std_logic := '0';
	signal sensor_we_shift :  std_logic := '0';
	signal sensor_we_valid :  std_logic := '0';

	signal cnt_fifo_in : std_logic_vector(15 downto 0);
	signal ack_fifo_in : std_logic;
	signal cnt_fifo_out  : std_logic_vector(15 downto 0);
	signal ack_fifo_out  : std_logic;

	-- puts
	signal fsm_mode	:  std_logic := '0';
	-- clock period definitions
	constant clk_period : time := 1 ns;

begin
	-- Instantiate the Unit Under Test (UUT)
	uut: fsm
	generic map (
			    NB_NEURONS => 1
		    )
	port map (
			 reset => reset,
			 clk => clk         ,
			 -- Control signals
			 ctrl_we_mode => ctrl_we_mode   ,
			 ctrl_we_shift => ctrl_we_shift  ,
			 ctrl_we_valid => ctrl_we_valid  ,
			 ctrl_accu_clear => ctrl_accu_clear,
			 ctrl_accu_add => ctrl_accu_add  ,
			 ctrl_shift_en => ctrl_shift_en  ,
			 ctrl_shift_copy => ctrl_shift_copy,
			 -- Address used for Read and Write
			 addr => addr           ,
			 -- Ports for Write Enable
			 n0_we_prev => n0_we_prev        ,
			 nN_we_next => nN_we_next        ,
			 -- Sensors, for synchronization with the controller
			 sensor_shift => sensor_shift   ,
			 sensor_copy => sensor_copy    ,
			 sensor_we_mode => sensor_we_mode ,
			 sensor_we_shift => sensor_we_shift,
			 sensor_we_valid => sensor_we_valid,
			 -- inputs
			 fsm_mode => fsm_mode,
			 -- in FIFO
			 cnt_fifo_in => cnt_fifo_in,
			 ack_fifo_in => ack_fifo_in,
			 cnt_fifo_out  => cnt_fifo_out,
			 ack_fifo_out  => ack_fifo_out
		 );       
	uut2: neuron
	port map (
			clk             => clk            ,
			-- Control signals
			ctrl_we_mode    => ctrl_we_mode   ,
			ctrl_we_shift   => ctrl_we_shift  ,
			ctrl_we_valid   => ctrl_we_valid  ,
			ctrl_accu_clear => ctrl_accu_clear,
			ctrl_accu_add   => ctrl_accu_add  ,
			ctrl_shift_en   => ctrl_shift_en  ,
			ctrl_shift_copy => ctrl_shift_copy,
			-- Address used for Read and Write
			addr            => addr           ,
			-- Ports for Write Enable
			we_prev         => n0_we_prev     ,
			we_next         => nN_we_next        ,
			write_data      => write_data     ,
			-- Data input, 2 bits
			data_in         => data_in        ,
			-- Scan chain to extract values
			sh_data_in      => sh_data_in     ,
			sh_data_out     => sh_data_out    ,
			-- Sensors, for synchronization with the controller
			sensor_shift    => sensor_shift   ,
			sensor_copy     => sensor_copy    ,
			sensor_we_mode  => sensor_we_mode ,
			sensor_we_shift => sensor_we_shift,
			sensor_we_valid => sensor_we_valid

		);


	-- Clock process definitions( clock with 50% duty cycle is generated here.
	clk_process :process
	begin
		clk <= '1';
		wait for clk_period/2;  --for 0.5 ns signal is '1'.
		clk <= '0';
		wait for clk_period/2;  --for next 0.5 ns signal is '0'.
	end process;

	----------------------
	-- Stimulus process --
	----------------------
	stim_proc: process
	begin         
		wait for 1 ns;
		
		-- reset component
		reset       <= '1';
		fsm_mode    <= '0';
		wait for clk_period;

		-- accu_mode
		reset       <= '0';
		fsm_mode    <= '1';
		sh_data_in <= X"00000000";
		wait for clk_period;
		write_data <= std_logic_vector(to_unsigned(1, write_data'length));
		sensor_we_valid <= '1';

		wait for 1000*clk_period;

		fsm_mode    <= '0';
		wait for clk_period;
		data_in <= std_logic_vector(to_unsigned(1, write_data'length));

		wait for 1000*clk_period;
		
	end process;

END;
