LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
USE ieee.std_logic_unsigned.all;
Library UNISIM;
use UNISIM.vcomponents.all;
library UNIMACRO;
use unimacro.Vcomponents.all;

-- entity declaration for your testbench.Dont declare any ports here
ENTITY test_bram IS 
	END test_bram;

ARCHITECTURE behavior OF test_bram IS
	SIGNAL do	: std_logic_vector(15 downto 0) ;
	SIGNAL addr	: std_logic_vector(9 downto 0) ; 
	SIGNAL di	: std_logic_vector(15 downto 0);
	SIGNAL en	: std_logic := '1';
	SIGNAL regce	: std_logic := '1';
	SIGNAL we	: std_logic_vector(1 downto 0) ;
	SIGNAL clk   : std_logic;
	SIGNAL rst   : std_logic;
   -- cLOCK PERIOD DEfinitions
	constant clk_period : time := 1 ns;
BEGIN
   -- Instantiate the Unit Under Test (UUT)
	uut: BRAM_SINGLE_MACRO 
	generic map (
			    BRAM_SIZE => "18Kb", -- Target BRAM, "18Kb" or "36Kb"
			    DEVICE => "7SERIES", -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
			    DO_REG => 0, -- Optional output register (0 or 1)
			    INIT => X"000000000000000000",   --  Initial values on output port
			    INIT_FILE => "NONE",
			    WRITE_WIDTH => 16,   -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
			    READ_WIDTH => 16,   -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
			    SRVAL => X"000000000000000000",   -- Set/Reset value for port output
			    WRITE_MODE => "WRITE_FIRST", -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
							 -- The following INIT_xx declarations specify the initial contents of the RAM
			    INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
			    INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
			    INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
			    INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
			    INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
			    INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
			    INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
			    INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
			    INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
			    INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
			    INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
			    INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
			    INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
			    INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
			    INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
			    INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
			    INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
			    INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
			    INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
			    INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
			    INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
			    INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
			    INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
			    INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
			    INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
			    INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
			    INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
			    INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
			    INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
			    INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
			    INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
			    INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
			    INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
			    INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
			    INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
			    INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
			    INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
			    INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
			    INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
			    INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
			    INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
			    INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
			    INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
			    INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
			    INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
			    INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
			    INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
			    INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
			    INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
			    INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
			    INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
			    INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
			    INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
			    INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
			    INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
			    INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
			    INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
			    INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
			    INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
			    INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
			    INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
			    INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
			    INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
			    INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000",
		    -- The next set of INIT_xx are valid when configured as 36Kb
			    INIT_40 => X"0000000000000000000000000000000000000000000000000000000000000000",
			    INIT_41 => X"0000000000000000000000000000000000000000000000000000000000000000",
			    INIT_42 => X"0000000000000000000000000000000000000000000000000000000000000000",
			    INIT_43 => X"0000000000000000000000000000000000000000000000000000000000000000",
			    INIT_44 => X"0000000000000000000000000000000000000000000000000000000000000000",
			    INIT_45 => X"0000000000000000000000000000000000000000000000000000000000000000",
			    INIT_46 => X"0000000000000000000000000000000000000000000000000000000000000000",
			    INIT_47 => X"0000000000000000000000000000000000000000000000000000000000000000",
			    INIT_48 => X"0000000000000000000000000000000000000000000000000000000000000000",
			    INIT_49 => X"0000000000000000000000000000000000000000000000000000000000000000",
			    INIT_4A => X"0000000000000000000000000000000000000000000000000000000000000000",
			    INIT_4B => X"0000000000000000000000000000000000000000000000000000000000000000",
			    INIT_4C => X"0000000000000000000000000000000000000000000000000000000000000000",
			    INIT_4D => X"0000000000000000000000000000000000000000000000000000000000000000",
			    INIT_4E => X"0000000000000000000000000000000000000000000000000000000000000000",
			    INIT_4F => X"0000000000000000000000000000000000000000000000000000000000000000",
			    INIT_50 => X"0000000000000000000000000000000000000000000000000000000000000000",
			    INIT_51 => X"0000000000000000000000000000000000000000000000000000000000000000",
			    INIT_52 => X"0000000000000000000000000000000000000000000000000000000000000000",
			    INIT_53 => X"0000000000000000000000000000000000000000000000000000000000000000",
			    INIT_54 => X"0000000000000000000000000000000000000000000000000000000000000000",
			    INIT_55 => X"0000000000000000000000000000000000000000000000000000000000000000",
			    INIT_56 => X"0000000000000000000000000000000000000000000000000000000000000000",
			    INIT_57 => X"0000000000000000000000000000000000000000000000000000000000000000",
			    INIT_58 => X"0000000000000000000000000000000000000000000000000000000000000000",
			    INIT_59 => X"0000000000000000000000000000000000000000000000000000000000000000",
			    INIT_5A => X"0000000000000000000000000000000000000000000000000000000000000000",
			    INIT_5B => X"0000000000000000000000000000000000000000000000000000000000000000",
			    INIT_5C => X"0000000000000000000000000000000000000000000000000000000000000000",
			    INIT_5D => X"0000000000000000000000000000000000000000000000000000000000000000",
			    INIT_5E => X"0000000000000000000000000000000000000000000000000000000000000000",
			    INIT_5F => X"0000000000000000000000000000000000000000000000000000000000000000",
			    INIT_60 => X"0000000000000000000000000000000000000000000000000000000000000000",
			    INIT_61 => X"0000000000000000000000000000000000000000000000000000000000000000",
			    INIT_62 => X"0000000000000000000000000000000000000000000000000000000000000000",
			    INIT_63 => X"0000000000000000000000000000000000000000000000000000000000000000",
			    INIT_64 => X"0000000000000000000000000000000000000000000000000000000000000000",
			    INIT_65 => X"0000000000000000000000000000000000000000000000000000000000000000",
			    INIT_66 => X"0000000000000000000000000000000000000000000000000000000000000000",
			    INIT_67 => X"0000000000000000000000000000000000000000000000000000000000000000",
			    INIT_68 => X"0000000000000000000000000000000000000000000000000000000000000000",
			    INIT_69 => X"0000000000000000000000000000000000000000000000000000000000000000",
			    INIT_6A => X"0000000000000000000000000000000000000000000000000000000000000000",
			    INIT_6B => X"0000000000000000000000000000000000000000000000000000000000000000",
			    INIT_6C => X"0000000000000000000000000000000000000000000000000000000000000000",
			    INIT_6D => X"0000000000000000000000000000000000000000000000000000000000000000",
			    INIT_6E => X"0000000000000000000000000000000000000000000000000000000000000000",
			    INIT_6F => X"0000000000000000000000000000000000000000000000000000000000000000",
			    INIT_70 => X"0000000000000000000000000000000000000000000000000000000000000000",
			    INIT_71 => X"0000000000000000000000000000000000000000000000000000000000000000",
			    INIT_72 => X"0000000000000000000000000000000000000000000000000000000000000000",
			    INIT_73 => X"0000000000000000000000000000000000000000000000000000000000000000",
			    INIT_74 => X"0000000000000000000000000000000000000000000000000000000000000000",
			    INIT_75 => X"0000000000000000000000000000000000000000000000000000000000000000",
			    INIT_76 => X"0000000000000000000000000000000000000000000000000000000000000000",
			    INIT_77 => X"0000000000000000000000000000000000000000000000000000000000000000",
			    INIT_78 => X"0000000000000000000000000000000000000000000000000000000000000000",
			    INIT_79 => X"0000000000000000000000000000000000000000000000000000000000000000",
			    INIT_7A => X"0000000000000000000000000000000000000000000000000000000000000000",
			    INIT_7B => X"0000000000000000000000000000000000000000000000000000000000000000",
			    INIT_7C => X"0000000000000000000000000000000000000000000000000000000000000000",
			    INIT_7D => X"0000000000000000000000000000000000000000000000000000000000000000",
			    INIT_7E => X"0000000000000000000000000000000000000000000000000000000000000000",
			    INIT_7F => X"0000000000000000000000000000000000000000000000000000000000000000",
		    -- The next set of INITP_xx are for the parity bits
			    INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
			    INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
			    INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
			    INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
			    INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
			    INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
			    INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
			    INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
		    -- The next set of INIT_xx are valid when configured as 36Kb
			    INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
			    INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
			    INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
			    INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
			    INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
			    INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
			    INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
			    INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000")
	port map (
			 DO => DO,      -- Output data, width defined by READ_WIDTH parameter
			 ADDR => ADDR,  -- Input address, width defined by read/write port depth
			 CLK => CLK,
			 DI => DI,
			 EN => EN,
			 REGCE => REGCE, -- 1-bit input output register enable
			 RST => RST,    -- 1-bit input reset
			 WE => WE       -- Input write enable, width defined by write port depth
		 );       

   -- Clock process definitions( clock with 50% duty cycle is generated here.
	clk_process :process
	begin
		clk <= '0';
		wait for clk_period/2;  --for 0.5 ns signal is '0'.
		clk <= '1';
		wait for clk_period/2;  --for next 0.5 ns signal is '1'.
	end process;
   -- Stimulus process
	stim_proc: process
	begin         
		wait for 1 ns;
		rst       <= '1';
		wait for 1 ns;
		rst       <= '0';

		wait for 1 ns;
		rst       <= '0';

		wait for 1 ns;
		rst       <= '0';

		wait for 1 ns;
		rst       <= '0';
		wait;
	end process;

END;
